// Copyright (C) Ganzin Technology - All Rights Reserved
// ---------------------------
// Unauthorized copying of this file, via any medium is strictly prohibited
// Proprietary and confidential
//
// Contributors
// ---------------------------
// En-Ho Shen <enhoshen@ganzin.com.tw>, [:VIM_EVAL:]strftime('%Y')[:END_EVAL:]

`ifndef __[:VIM_EVAL:]toupper(''.expand("<afile>:t:r"))[:END_EVAL:]_SV__
`define __[:VIM_EVAL:]toupper(''.expand("<afile>:t:r"))[:END_EVAL:]_SV__

// packages

// sub-modules

`endif //__[:VIM_EVAL:]toupper(''.expand("<afile>:t:r"))[:END_EVAL:]_SV__
