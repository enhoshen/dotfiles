// packages

// sub-modules

module [:VIM_EVAL:]''.expand("<afile>:r")[:END_EVAL:]
#(
)(
     input i_clk
    ,input i_rst_n
);
    //====================
    //     parameter 
    //====================
    //====================
    //       logic 
    //====================
    //====================
    //   combinational 
    //====================
    //====================
    //     sequential 
    //====================

endmodule
